**.subckt INV_tb
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
Vdd Vdd 0 3.3
Vin Vin 0 dc pulse(0 3.3 0 1p 1p 100p 200p)
X1 Vdd Vout Vin 0 INV


.temp -40
.options tnom=-40


.control
tran 1p 400p
meas tran tphl TRIG v(Vin) VAL={0.5*3.3} RISE=2 TARG v(Vout) VAL={0.5*3.3} FALL=2
meas tran tplh TRIG v(Vin) VAL={0.5*3.3} FALL=1 TARG v(Vout) VAL={0.5*3.3} RISE=1
print {(tplh+tphl)/2}
wrdata ../run_smoke_2023-11-25_14:51:02.640025/simulation/inv_W0.22_L0.28_T-40_ff.csv {(tplh+tphl)/2}
.endc


.include "../../design.ngspice"
.lib "../../sm141064.ngspice" ff


.subckt INV  VDD Vout Vin GND
XM1 Vout Vin GND GND nmos_3p3 W=0.22u L=0.28u
*ad=p pd=u as=p ps=u
XM2 Vout Vin VDD VDD pmos_3p3 W = 0.33u L = 0.28u
*ad=u pd=u as=u ps=u
.ends

.end